library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

entity calc is
port(
    clk : in std_logic;
    reset : in std_logic
);
end entity;

architecture rtl of calc is
begin

process(all) begin
  if rising_edge(clk) then
  end if;
end process;

end architecture;

